LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE work.aes_pack.ALL;
ENTITY mixcolumn IS
	PORT(
		a 	: IN  std_logic_vector(127 DOWNTO 0);
		mcl : OUT std_logic_vector(127 DOWNTO 0)
	);
END mixcolumn;
ARCHITECTURE dataflow OF mixcolumn IS
BEGIN
	mcl(127 DOWNTO 120) <= mcl32(a(127 DOWNTO 120),a(119 DOWNTO 112),a(111 DOWNTO 104),a(103 DOWNTO 96));
	mcl(119 DOWNTO 112) <= mcl32(a(119 DOWNTO 112),a(111 DOWNTO 104),a(103 DOWNTO 96),a(127 DOWNTO 120));
	mcl(111 DOWNTO 104) <= mcl32(a(111 DOWNTO 104),a(103 DOWNTO 96),a(127 DOWNTO 120),a(119 DOWNTO 112));
	mcl(103 DOWNTO 96)  <= mcl32(a(103 DOWNTO 96),a(127 DOWNTO 120),a(119 DOWNTO 112),a(111 DOWNTO 104));
	mcl(95  DOWNTO 88)  <= mcl32(a(95 DOWNTO 88),a(87 DOWNTO 80),a(79 DOWNTO 72),a(71 DOWNTO 64));
	mcl(87  DOWNTO 80)  <= mcl32(a(87 DOWNTO 80),a(79 DOWNTO 72),a(71 DOWNTO 64),a(95 DOWNTO 88));
	mcl(79  DOWNTO 72)  <= mcl32(a(79 DOWNTO 72),a(71 DOWNTO 64),a(95 DOWNTO 88),a(87 DOWNTO 80));
	mcl(71  DOWNTO 64)  <= mcl32(a(71 DOWNTO 64),a(95 DOWNTO 88),a(87 DOWNTO 80),a(79 DOWNTO 72));
	mcl(63  DOWNTO 56)  <= mcl32(a(63 DOWNTO 56),a(55 DOWNTO 48),a(47 DOWNTO 40),a(39 DOWNTO 32));
	mcl(55  DOWNTO 48)  <= mcl32(a(55 DOWNTO 48),a(47 DOWNTO 40),a(39 DOWNTO 32),a(63 DOWNTO 56));
	mcl(47  DOWNTO 40)  <= mcl32(a(47 DOWNTO 40),a(39 DOWNTO 32),a(63 DOWNTO 56),a(55 DOWNTO 48));
	mcl(39  DOWNTO 32)  <= mcl32(a(39 DOWNTO 32),a(63 DOWNTO 56),a(55 DOWNTO 48),a(47 DOWNTO 40));
	mcl(31  DOWNTO 24)  <= mcl32(a(31 DOWNTO 24),a(23 DOWNTO 16),a(15 DOWNTO 8),a(7 DOWNTO 0));
	mcl(23  DOWNTO 16)  <= mcl32(a(23 DOWNTO 16),a(15 DOWNTO 8),a(7 DOWNTO 0),a(31 DOWNTO 24));
	mcl(15  DOWNTO 8)   <= mcl32(a(15 DOWNTO 8),a(7 DOWNTO 0),a(31 DOWNTO 24),a(23 DOWNTO 16));
	mcl(7   DOWNTO 0)   <= mcl32(a(7 DOWNTO 0),a(31 DOWNTO 24),a(23 DOWNTO 16),a(15 DOWNTO 8));
END dataflow;