LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE work.aes_pack.ALL;
ENTITY sbox IS
	PORT(
		a 	: IN  std_logic_vector(7 DOWNTO 0);
		c 	: OUT std_logic_vector(7 DOWNTO 0)
	);
END sbox;
ARCHITECTURE behavioral OF sbox IS
BEGIN 
	PROCESS(a)
	BEGIN
		CASE a IS
			WHEN X"00" 	=> c <= X"63";
			WHEN X"01" 	=> c <= X"7c";
			WHEN X"02" 	=> c <= X"77";
			WHEN X"03" 	=> c <= X"7b";
			WHEN X"04" 	=> c <= X"f2";
			WHEN X"05" 	=> c <= X"6b";
			WHEN X"06" 	=> c <= X"6f";
			WHEN X"07" 	=> c <= X"c5";
			WHEN X"08" 	=> c <= X"30";
			WHEN X"09" 	=> c <= X"01";
			WHEN X"0a" 	=> c <= X"67";
			WHEN X"0b" 	=> c <= X"2b";
			WHEN X"0c" 	=> c <= X"fe";
			WHEN X"0d" 	=> c <= X"d7";
			WHEN X"0e" 	=> c <= X"ab";
			WHEN X"0f" 	=> c <= X"76";
			WHEN X"10" 	=> c <= X"ca";
			WHEN X"11" 	=> c <= X"82";
			WHEN X"12" 	=> c <= X"c9";
			WHEN X"13" 	=> c <= X"7d";
			WHEN X"14" 	=> c <= X"fa";
			WHEN X"15" 	=> c <= X"59";
			WHEN X"16" 	=> c <= X"47";
			WHEN X"17" 	=> c <= X"f0";
			WHEN X"18" 	=> c <= X"ad";
			WHEN X"19" 	=> c <= X"d4";
			WHEN X"1a" 	=> c <= X"a2";
			WHEN X"1b" 	=> c <= X"af";
			WHEN X"1c" 	=> c <= X"9c";
			WHEN X"1d" 	=> c <= X"a4";
			WHEN X"1e" 	=> c <= X"72";
			WHEN X"1f" 	=> c <= X"c0";
			WHEN X"20" 	=> c <= X"b7";
			WHEN X"21" 	=> c <= X"fd";
			WHEN X"22" 	=> c <= X"93";
			WHEN X"23" 	=> c <= X"26";
			WHEN X"24" 	=> c <= X"36";
			WHEN X"25" 	=> c <= X"3f";
			WHEN X"26" 	=> c <= X"f7";
			WHEN X"27" 	=> c <= X"cc";
			WHEN X"28" 	=> c <= X"34";
			WHEN X"29" 	=> c <= X"a5";
			WHEN X"2a" 	=> c <= X"e5";
			WHEN X"2b" 	=> c <= X"f1";
			WHEN X"2c" 	=> c <= X"71";
			WHEN X"2d" 	=> c <= X"d8";
			WHEN X"2e" 	=> c <= X"31";
			WHEN X"2f" 	=> c <= X"15";
			WHEN X"30" 	=> c <= X"04";
			WHEN X"31" 	=> c <= X"c7";
			WHEN X"32" 	=> c <= X"23";
			WHEN X"33" 	=> c <= X"c3";
			WHEN X"34" 	=> c <= X"18";
			WHEN X"35" 	=> c <= X"96";
			WHEN X"36" 	=> c <= X"05";
			WHEN X"37" 	=> c <= X"9a";
			WHEN X"38" 	=> c <= X"07";
			WHEN X"39" 	=> c <= X"12";
			WHEN X"3a" 	=> c <= X"80";
			WHEN X"3b" 	=> c <= X"e2";
			WHEN X"3c" 	=> c <= X"eb";
			WHEN X"3d" 	=> c <= X"27";
			WHEN X"3e" 	=> c <= X"b2";
			WHEN X"3f" 	=> c <= X"75";
			WHEN X"40" 	=> c <= X"09";
			WHEN X"41" 	=> c <= X"83";
			WHEN X"42" 	=> c <= X"2c";
			WHEN X"43" 	=> c <= X"1a";
			WHEN X"44" 	=> c <= X"1b";
			WHEN X"45" 	=> c <= X"6e";
			WHEN X"46" 	=> c <= X"5a";
			WHEN X"47" 	=> c <= X"a0";
			WHEN X"48" 	=> c <= X"52";
			WHEN X"49" 	=> c <= X"3b";
			WHEN X"4a" 	=> c <= X"d6";
			WHEN X"4b" 	=> c <= X"b3";
			WHEN X"4c" 	=> c <= X"29";
			WHEN X"4d" 	=> c <= X"e3";
			WHEN X"4e" 	=> c <= X"2f";
			WHEN X"4f" 	=> c <= X"84";
			WHEN X"50" 	=> c <= X"53";
			WHEN X"51" 	=> c <= X"d1";
			WHEN X"52" 	=> c <= X"00";
			WHEN X"53" 	=> c <= X"ed";
			WHEN X"54" 	=> c <= X"20";
			WHEN X"55" 	=> c <= X"fc";
			WHEN X"56" 	=> c <= X"b1";
			WHEN X"57" 	=> c <= X"5b";
			WHEN X"58" 	=> c <= X"6a";
			WHEN X"59" 	=> c <= X"cb";
			WHEN X"5a" 	=> c <= X"be";
			WHEN X"5b" 	=> c <= X"39";
			WHEN X"5c" 	=> c <= X"4a";
			WHEN X"5d" 	=> c <= X"4c";
			WHEN X"5e" 	=> c <= X"58";
			WHEN X"5f" 	=> c <= X"cf";
			WHEN X"60" 	=> c <= X"d0";
			WHEN X"61" 	=> c <= X"ef";
			WHEN X"62" 	=> c <= X"aa";
			WHEN X"63" 	=> c <= X"fb";
			WHEN X"64" 	=> c <= X"43";
			WHEN X"65" 	=> c <= X"4d";
			WHEN X"66" 	=> c <= X"33";
			WHEN X"67" 	=> c <= X"85";
			WHEN X"68" 	=> c <= X"45";
			WHEN X"69" 	=> c <= X"f9";
			WHEN X"6a" 	=> c <= X"02";
			WHEN X"6b" 	=> c <= X"7f";
			WHEN X"6c" 	=> c <= X"50";
			WHEN X"6d" 	=> c <= X"3c";
			WHEN X"6e" 	=> c <= X"9f";
			WHEN X"6f" 	=> c <= X"a8";
			WHEN X"70" 	=> c <= X"51";
			WHEN X"71" 	=> c <= X"a3";
			WHEN X"72" 	=> c <= X"40";
			WHEN X"73" 	=> c <= X"8f";
			WHEN X"74" 	=> c <= X"92";
			WHEN X"75" 	=> c <= X"9d";
			WHEN X"76" 	=> c <= X"38";
			WHEN X"77" 	=> c <= X"f5";
			WHEN X"78" 	=> c <= X"bc";
			WHEN X"79" 	=> c <= X"b6";
			WHEN X"7a" 	=> c <= X"da";
			WHEN X"7b" 	=> c <= X"21";
			WHEN X"7c" 	=> c <= X"10";
			WHEN X"7d" 	=> c <= X"ff";
			WHEN X"7e" 	=> c <= X"f3";
			WHEN X"7f" 	=> c <= X"d2";
			WHEN X"80" 	=> c <= X"cd";
			WHEN X"81" 	=> c <= X"0c";
			WHEN X"82" 	=> c <= X"13";
			WHEN X"83" 	=> c <= X"ec";
			WHEN X"84" 	=> c <= X"5f";
			WHEN X"85" 	=> c <= X"97";
			WHEN X"86" 	=> c <= X"44";
			WHEN X"87" 	=> c <= X"17";
			WHEN X"88" 	=> c <= X"c4";
			WHEN X"89" 	=> c <= X"a7";
			WHEN X"8a" 	=> c <= X"7e";
			WHEN X"8b" 	=> c <= X"3d";
			WHEN X"8c" 	=> c <= X"64";
			WHEN X"8d" 	=> c <= X"5d";
			WHEN X"8e" 	=> c <= X"19";
			WHEN X"8f" 	=> c <= X"73";
			WHEN X"90" 	=> c <= X"60";
			WHEN X"91" 	=> c <= X"81";
			WHEN X"92" 	=> c <= X"4f";
			WHEN X"93" 	=> c <= X"dc";
			WHEN X"94" 	=> c <= X"22";
			WHEN X"95" 	=> c <= X"2a";
			WHEN X"96" 	=> c <= X"90";
			WHEN X"97" 	=> c <= X"88";
			WHEN X"98" 	=> c <= X"46";
			WHEN X"99" 	=> c <= X"ee";
			WHEN X"9a" 	=> c <= X"b8";
			WHEN X"9b" 	=> c <= X"14";
			WHEN X"9c" 	=> c <= X"de";
			WHEN X"9d" 	=> c <= X"5e";
			WHEN X"9e" 	=> c <= X"0b";
			WHEN X"9f" 	=> c <= X"db";
			WHEN X"a0" 	=> c <= X"e0";
			WHEN X"a1" 	=> c <= X"32";
			WHEN X"a2" 	=> c <= X"3a";
			WHEN X"a3" 	=> c <= X"0a";
			WHEN X"a4" 	=> c <= X"49";
			WHEN X"a5" 	=> c <= X"06";
			WHEN X"a6" 	=> c <= X"24";
			WHEN X"a7" 	=> c <= X"5c";
			WHEN X"a8" 	=> c <= X"c2";
			WHEN X"a9" 	=> c <= X"d3";
			WHEN X"aa" 	=> c <= X"ac";
			WHEN X"ab" 	=> c <= X"62";
			WHEN X"ac" 	=> c <= X"91";
			WHEN X"ad" 	=> c <= X"95";
			WHEN X"ae" 	=> c <= X"e4";
			WHEN X"af" 	=> c <= X"79";
			WHEN X"b0" 	=> c <= X"e7";
			WHEN X"b1" 	=> c <= X"c8";
			WHEN X"b2" 	=> c <= X"37";
			WHEN X"b3" 	=> c <= X"6d";
			WHEN X"b4" 	=> c <= X"8d";
			WHEN X"b5" 	=> c <= X"d5";
			WHEN X"b6" 	=> c <= X"4e";
			WHEN X"b7" 	=> c <= X"a9";
			WHEN X"b8" 	=> c <= X"6c";
			WHEN X"b9" 	=> c <= X"56";
			WHEN X"ba" 	=> c <= X"f4";
			WHEN X"bb" 	=> c <= X"ea";
			WHEN X"bc" 	=> c <= X"65";
			WHEN X"bd" 	=> c <= X"7a";
			WHEN X"be" 	=> c <= X"ae";
			WHEN X"bf" 	=> c <= X"08";
			WHEN X"c0" 	=> c <= X"ba";
			WHEN X"c1" 	=> c <= X"78";
			WHEN X"c2" 	=> c <= X"25";
			WHEN X"c3" 	=> c <= X"2e";
			WHEN X"c4" 	=> c <= X"1c";
			WHEN X"c5" 	=> c <= X"a6";
			WHEN X"c6" 	=> c <= X"b4";
			WHEN X"c7" 	=> c <= X"c6";
			WHEN X"c8" 	=> c <= X"e8";
			WHEN X"c9" 	=> c <= X"dd";
			WHEN X"ca" 	=> c <= X"74";
			WHEN X"cb" 	=> c <= X"1f";
			WHEN X"cc" 	=> c <= X"4b";
			WHEN X"cd" 	=> c <= X"bd";
			WHEN X"ce" 	=> c <= X"8b";
			WHEN X"cf" 	=> c <= X"8a";
			WHEN X"d0" 	=> c <= X"70";
			WHEN X"d1" 	=> c <= X"3e";
			WHEN X"d2" 	=> c <= X"b5";
			WHEN X"d3" 	=> c <= X"66";
			WHEN X"d4" 	=> c <= X"48";
			WHEN X"d5" 	=> c <= X"03";
			WHEN X"d6" 	=> c <= X"f6";
			WHEN X"d7" 	=> c <= X"0e";
			WHEN X"d8" 	=> c <= X"61";
			WHEN X"d9" 	=> c <= X"35";
			WHEN X"da" 	=> c <= X"57";
			WHEN X"db" 	=> c <= X"b9";
			WHEN X"dc" 	=> c <= X"86";
			WHEN X"dd" 	=> c <= X"c1";
			WHEN X"de" 	=> c <= X"1d";
			WHEN X"df" 	=> c <= X"9e";
			WHEN X"e0" 	=> c <= X"e1";
			WHEN X"e1" 	=> c <= X"f8";
			WHEN X"e2" 	=> c <= X"98";
			WHEN X"e3" 	=> c <= X"11";
			WHEN X"e4" 	=> c <= X"69";
			WHEN X"e5" 	=> c <= X"d9";
			WHEN X"e6" 	=> c <= X"8e";
			WHEN X"e7" 	=> c <= X"94";
			WHEN X"e8" 	=> c <= X"9b";
			WHEN X"e9" 	=> c <= X"1e";
			WHEN X"ea" 	=> c <= X"87";
			WHEN X"eb" 	=> c <= X"e9";
			WHEN X"ec" 	=> c <= X"ce";
			WHEN X"ed" 	=> c <= X"55";
			WHEN X"ee" 	=> c <= X"28";
			WHEN X"ef" 	=> c <= X"df";
			WHEN X"f0" 	=> c <= X"8c";
			WHEN X"f1" 	=> c <= X"a1";
			WHEN X"f2" 	=> c <= X"89";
			WHEN X"f3" 	=> c <= X"0d";
			WHEN X"f4" 	=> c <= X"bf";
			WHEN X"f5" 	=> c <= X"e6";
			WHEN X"f6" 	=> c <= X"42";
			WHEN X"f7" 	=> c <= X"68";
			WHEN X"f8" 	=> c <= X"41";
			WHEN X"f9" 	=> c <= X"99";
			WHEN X"fa" 	=> c <= X"2d";
			WHEN X"fb" 	=> c <= X"0f";
			WHEN X"fc" 	=> c <= X"b0";
			WHEN X"fd" 	=> c <= X"54";
			WHEN X"fe" 	=> c <= X"bb";
			WHEN OTHERS => c <= X"16";
		END CASE;
	END PROCESS;
END behavioral;